module point_doubling ();

endmodule // point_doubling
