module point_addition ();

endmodule // point_addition
